library verilog;
use verilog.vl_types.all;
entity portao_vlg_vec_tst is
end portao_vlg_vec_tst;
